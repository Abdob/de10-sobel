module SOBEL(GRAY,OUTPUT); 

input [7:0] GRAY;

output [7:0] OUTPUT; 
 
assign OUTPUT = GRAY;

endmodule